* Qucs 0.0.22 /usr/share/qucs-s/examples/ngspice/BJT.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.22  /usr/share/qucs-s/examples/ngspice/BJT.sch
.PARAM Rload=47k
Q2N2222A_1 _net1 _net0 _net2 QMOD_Q2N2222A_1 AREA=1 TEMP=26.85
.MODEL QMOD_Q2N2222A_1 npn (Is=8.11e-14 Nf=1 Nr=1 Ikf=0.5 Ikr=0.225 Vaf=113 Var=24 Ise=1.06e-11 Ne=2 Isc=0 Nc=2 Bf=205 Br=4 Rbm=0 Irb=0 Rc=0.137 Re=0.343 Rb=1.37 Cje=2.95e-11 Vje=0.75 Mje=0.33 Cjc=1.52e-11 Vjc=0.75 Mjc=0.33 Xcjc=1 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=3.97e-10 Xtf=0 Vtf=0 Itf=0 Tr=8.5e-08 Kf=0 Af=1 Ptf=0 Xtb=1.5 Xti=3 Eg=1.11 Tnom=26.85 )
R1 0 _net0  2K
R2 0 _net2  470
C1 in _net0  0.1U 
R3 _net0 _net3  24K
C2 _net1 out  0.1U 
V1 _net4 0 DC 12
R5 _net1 _net3  4.7K
V2 in 0 DC 0 SIN(0 200M 4K 0 0 0) AC 200M
R4 0 out  {RLOAD}
VPr1 _net4 _net3 DC 0
.control
*echo "" > spice4qucs.cir.noise
*echo "" > spice4qucs.cir.pz
set gnuplot_terminal=png

let Rload=47k
tran 1e-06 0.001 0 
let Pwr=(V(out)*V(out))/Rload
write circuits/qucs-npn-tran.data VPr1#branch v(in) v(out) Pwr
gnuplot circuits/qucs-npn-pwr Pwr
gnuplot circuits/qucs-npn-voltage v(in) v(out)
destroy all
reset

let Rload=47k
ac dec 21 100 10meg 
let K=V(out)/V(in)
write circuits/qucs-npn-ac.data VPr1#branch v(in) v(out)  K
gnuplot circuits/qucs-npn-gain v(in) v(out) K
destroy all
reset

exit
.endc
.END
